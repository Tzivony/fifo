package fifo_pack;
	typedef enum {
		CNTR,
		CALC,
		NONE
	} fl_type_e;
	
endpackage : fifo_pack